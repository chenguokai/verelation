module SRAMTemplate(
endmodule
